module main

import log4v

// TODO: add log4v benchmark in a multi-threaded console app ... wip

fn main() {
}
