module main

import log4v

// TODO: add log4v benchmark in a console app ...

fn main() {
}
